library ieee;
use ieee.std_logic_1164.all;


entity Diviseur_frequence is   port( 
	clkin : in std_logic;
	clkout : out std_logic);
end Diviseur_frequence ;